module Game_End(
    input            vga_clk_25,      
    input            rst_n,             
    input     [ 9:0] pixel_xpos,        
    input     [ 9:0] pixel_ypos,       
    input     [ 5:0] game_score,        
    
    output reg[15:0] pixel_data       
);
 

parameter   H_DISP = 10'd640;           
parameter   V_DISP = 10'd480;           

localparam  ROW1_X  = 10'd250;          
localparam  ROW1_Y  = 10'd180;          
localparam  ROW1_H  = 10'd160;          
localparam  ROW1_V  = 10'd32;           

localparam  ROW2_X  = 10'd280;          
localparam  ROW2_Y  = 10'd230;          
localparam  ROW2_H  = 10'd48;           
localparam  ROW2_V  = 10'd16;           

localparam  ROW3_X  = 10'd340;          
localparam  ROW3_Y  = 10'd230;          
localparam  ROW3_H  = 10'd16;           
localparam  ROW3_V  = 10'd16;           

localparam  WHITE  = 16'hFFFF;  
localparam  BLANK  = 16'h0000;  
localparam  RED    = 16'hF800;  
localparam  GREEN  = 16'h0400;  
localparam  BLUE   = 16'h001F;  
localparam  YELLOW = 16'hFFE0;  
localparam  PURPLE = 16'h8010;  
localparam  BROWN  = 16'hE618;  

reg [159:0] row_1 [31:0];   
reg [ 47:0] row_2 [15:0];   
reg [ 15:0] row_3 [15:0];   

wire [9:0] x1_cnt;          
wire [9:0] y1_cnt;          
wire [9:0] x2_cnt;          
wire [9:0] y2_cnt;          
wire [9:0] x3_cnt;          
wire [9:0] y3_cnt;          


 

assign x1_cnt = pixel_xpos - ROW1_X;
assign y1_cnt = pixel_ypos - ROW1_Y;
assign x2_cnt = pixel_xpos - ROW2_X;
assign y2_cnt = pixel_ypos - ROW2_Y;
assign x3_cnt = pixel_xpos - ROW3_X;
assign y3_cnt = pixel_ypos - ROW3_Y;


always @(posedge vga_clk_25)
begin
    row_1[0]  <= 160'h0000000000000000000000000000000000000000;
    row_1[1]  <= 160'h0000000000000000000000000000000000000000;
    row_1[2]  <= 160'h0000000000000000000000000000000000000000;
    row_1[3]  <= 160'h0000000000000000000000000000000000000000;
    row_1[4]  <= 160'h0000000000000000000000000000000000000000;
    row_1[5]  <= 160'h0000000000000000000000000000000000000000;
    row_1[6]  <= 160'h03C00380F00F7FFC0000000003C07C1E7FFC7FE0;
    row_1[7]  <= 160'h0C300380381C180C000000000C30180C180C1838;
    row_1[8]  <= 160'h08100380381C1804000000001818180818041818;
    row_1[9]  <= 160'h18180380381C180200000000100818081802180C;
    row_1[10] <= 160'h300804C0381C180200000000300C18081802180C;
    row_1[11] <= 160'h300804C0382C180000000000300C0C101800180C;
    row_1[12] <= 160'h200004C02C2C18000000000060040C101800180C;
    row_1[13] <= 160'h600004C02C2C18100000000060060C101810180C;
    row_1[14] <= 160'h60000C402C2C18100000000060060C1018101818;
    row_1[15] <= 160'h600008602C4C18300000000060060C2018301830;
    row_1[16] <= 160'h600008602C4C1FF000000000600606201FF01FE0;
    row_1[17] <= 160'h60000860264C18300000000060060620183018C0;
    row_1[18] <= 160'h607E1820264C18100000000060060620181018C0;
    row_1[19] <= 160'h60181FF0264C1810000000006006064018101860;
    row_1[20] <= 160'h60181030268C1800000000006006034018001860;
    row_1[21] <= 160'h20181030228C1800000000002006034018001860;
    row_1[22] <= 160'h30181030238C180000000000300C034018001830;
    row_1[23] <= 160'h30182018238C180200000000300C038018021830;
    row_1[24] <= 160'h10182018230C1802000000001008018018021830;
    row_1[25] <= 160'h18182018230C1804000000001818018018041818;
    row_1[26] <= 160'h0C20601C210C180C000000000C300100180C1818;
    row_1[27] <= 160'h07C0F83EF13F7FFC0000000003C001007FFC7E1E;
    row_1[28] <= 160'h0000000000000000000000000000000000000000;
    row_1[29] <= 160'h0000000000000000000000000000000000000000;
    row_1[30] <= 160'h0000000000000000000000000000000000000000;
    row_1[31] <= 160'h0000000000000000000000000000000000000000;
    
    row_2[0]  <= 48'h000000000000;
    row_2[1]  <= 48'h000000000000;
    row_2[2]  <= 48'h000000000000;
    row_2[3]  <= 48'h3E3E38FCFC00;
    row_2[4]  <= 48'h424244424200;
    row_2[5]  <= 48'h424282424800;
    row_2[6]  <= 48'h408082424818;
    row_2[7]  <= 48'h2080827C7818;
    row_2[8]  <= 48'h188082484800;
    row_2[9]  <= 48'h048082484800;
    row_2[10] <= 48'h028082444000;
    row_2[11] <= 48'h424282444200;
    row_2[12] <= 48'h424444424318;
    row_2[13] <= 48'h7C3838E3FC18;
    row_2[14] <= 48'h000000000000;
    row_2[15] <= 48'h000000000000;
    
    case(game_score)
        6'd0:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h1818;
            row_3[4]  <= 16'h2424;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4242;  row_3[7]  <= 16'h4242;
            row_3[8]  <= 16'h4242;  row_3[9]  <= 16'h4242;  row_3[10] <= 16'h4242;  row_3[11] <= 16'h4242;
            row_3[12] <= 16'h2424;  row_3[13] <= 16'h1818;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd1:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h1808;
            row_3[4]  <= 16'h2438;  row_3[5]  <= 16'h4208;  row_3[6]  <= 16'h4208;  row_3[7]  <= 16'h4208;
            row_3[8]  <= 16'h4208;  row_3[9]  <= 16'h4208;  row_3[10] <= 16'h4208;  row_3[11] <= 16'h4208;
            row_3[12] <= 16'h2408;  row_3[13] <= 16'h183E;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd2:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h183C;
            row_3[4]  <= 16'h2442;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4242;  row_3[7]  <= 16'h4202;
            row_3[8]  <= 16'h4204;  row_3[9]  <= 16'h4208;  row_3[10] <= 16'h4210;  row_3[11] <= 16'h4220;
            row_3[12] <= 16'h2442;  row_3[13] <= 16'h187E;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd3:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h183C;
            row_3[4]  <= 16'h2442;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4202;  row_3[7]  <= 16'h4204;
            row_3[8]  <= 16'h4218;  row_3[9]  <= 16'h4204;  row_3[10] <= 16'h4202;  row_3[11] <= 16'h4242;
            row_3[12] <= 16'h2442;  row_3[13] <= 16'h183C;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd4:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h1804;
            row_3[4]  <= 16'h240C;  row_3[5]  <= 16'h420C;  row_3[6]  <= 16'h4214;  row_3[7]  <= 16'h4224;
            row_3[8]  <= 16'h4224;  row_3[9]  <= 16'h4244;  row_3[10] <= 16'h427F;  row_3[11] <= 16'h4204;
            row_3[12] <= 16'h2404;  row_3[13] <= 16'h181F;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd5:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h187E;
            row_3[4]  <= 16'h2440;  row_3[5]  <= 16'h4240;  row_3[6]  <= 16'h4240;  row_3[7]  <= 16'h4278;
            row_3[8]  <= 16'h4244;  row_3[9]  <= 16'h4202;  row_3[10] <= 16'h4202;  row_3[11] <= 16'h4242;
            row_3[12] <= 16'h2444;  row_3[13] <= 16'h1838;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd6:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h1818;
            row_3[4]  <= 16'h2424;  row_3[5]  <= 16'h4240;  row_3[6]  <= 16'h4240;  row_3[7]  <= 16'h425C;
            row_3[8]  <= 16'h4262;  row_3[9]  <= 16'h4242;  row_3[10] <= 16'h4242;  row_3[11] <= 16'h4242;
            row_3[12] <= 16'h2422;  row_3[13] <= 16'h181C;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd7:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h187E;
            row_3[4]  <= 16'h2442;  row_3[5]  <= 16'h4204;  row_3[6]  <= 16'h4204;  row_3[7]  <= 16'h4208;
            row_3[8]  <= 16'h4208;  row_3[9]  <= 16'h4210;  row_3[10] <= 16'h4210;  row_3[11] <= 16'h4210;
            row_3[12] <= 16'h2410;  row_3[13] <= 16'h1810;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd8:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h183C;
            row_3[4]  <= 16'h2442;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4242;  row_3[7]  <= 16'h4224;
            row_3[8]  <= 16'h4218;  row_3[9]  <= 16'h4224;  row_3[10] <= 16'h4242;  row_3[11] <= 16'h4242;
            row_3[12] <= 16'h2442;  row_3[13] <= 16'h183C;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd9:  begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h1838;
            row_3[4]  <= 16'h2444;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4242;  row_3[7]  <= 16'h4242;
            row_3[8]  <= 16'h4246;  row_3[9]  <= 16'h423A;  row_3[10] <= 16'h4202;  row_3[11] <= 16'h4202;
            row_3[12] <= 16'h2424;  row_3[13] <= 16'h1818;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd10: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h0818;
            row_3[4]  <= 16'h3824;  row_3[5]  <= 16'h0842;  row_3[6]  <= 16'h0842;  row_3[7]  <= 16'h0842;
            row_3[8]  <= 16'h0842;  row_3[9]  <= 16'h0842;  row_3[10] <= 16'h0842;  row_3[11] <= 16'h0842;
            row_3[12] <= 16'h0842;  row_3[13] <= 16'h3E18;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd11: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h0808;
            row_3[4]  <= 16'h3838;  row_3[5]  <= 16'h0808;  row_3[6]  <= 16'h0808;  row_3[7]  <= 16'h0808;
            row_3[8]  <= 16'h0808;  row_3[9]  <= 16'h0808;  row_3[10] <= 16'h0808;  row_3[11] <= 16'h0808;
            row_3[12] <= 16'h0808;  row_3[13] <= 16'h3E3E;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd12: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h083C;
            row_3[4]  <= 16'h3842;  row_3[5]  <= 16'h0842;  row_3[6]  <= 16'h0842;  row_3[7]  <= 16'h0802;
            row_3[8]  <= 16'h0804;  row_3[9]  <= 16'h0808;  row_3[10] <= 16'h0810;  row_3[11] <= 16'h0820;
            row_3[12] <= 16'h0842;  row_3[13] <= 16'h3E7E;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd13: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h083C;
            row_3[4]  <= 16'h3842;  row_3[5]  <= 16'h0842;  row_3[6]  <= 16'h0802;  row_3[7]  <= 16'h0804;
            row_3[8]  <= 16'h0818;  row_3[9]  <= 16'h0804;  row_3[10] <= 16'h0802;  row_3[11] <= 16'h0842;
            row_3[12] <= 16'h0842;  row_3[13] <= 16'h3E3C;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd14: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h0804;
            row_3[4]  <= 16'h380C;  row_3[5]  <= 16'h080C;  row_3[6]  <= 16'h0814;  row_3[7]  <= 16'h0824;
            row_3[8]  <= 16'h0824;  row_3[9]  <= 16'h0844;  row_3[10] <= 16'h087F;  row_3[11] <= 16'h0804;
            row_3[12] <= 16'h0804;  row_3[13] <= 16'h3E1F;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd15: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h087E;
            row_3[4]  <= 16'h3840;  row_3[5]  <= 16'h0840;  row_3[6]  <= 16'h0840;  row_3[7]  <= 16'h0878;
            row_3[8]  <= 16'h0844;  row_3[9]  <= 16'h0802;  row_3[10] <= 16'h0802;  row_3[11] <= 16'h0842;
            row_3[12] <= 16'h0844;  row_3[13] <= 16'h3E38;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd16: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h0818;
            row_3[4]  <= 16'h3824;  row_3[5]  <= 16'h0840;  row_3[6]  <= 16'h0840;  row_3[7]  <= 16'h085C;
            row_3[8]  <= 16'h0862;  row_3[9]  <= 16'h0842;  row_3[10] <= 16'h0842;  row_3[11] <= 16'h0842;
            row_3[12] <= 16'h0822;  row_3[13] <= 16'h3E1C;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd17: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h087E;
            row_3[4]  <= 16'h3842;  row_3[5]  <= 16'h0804;  row_3[6]  <= 16'h0804;  row_3[7]  <= 16'h0808;
            row_3[8]  <= 16'h0808;  row_3[9]  <= 16'h0810;  row_3[10] <= 16'h0810;  row_3[11] <= 16'h0810;
            row_3[12] <= 16'h0810;  row_3[13] <= 16'h3E10;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd18: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h083C;
            row_3[4]  <= 16'h3842;  row_3[5]  <= 16'h0842;  row_3[6]  <= 16'h0842;  row_3[7]  <= 16'h0824;
            row_3[8]  <= 16'h0818;  row_3[9]  <= 16'h0824;  row_3[10] <= 16'h0842;  row_3[11] <= 16'h0842;
            row_3[12] <= 16'h0842;  row_3[13] <= 16'h3E3C;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd19: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h0838;
            row_3[4]  <= 16'h3844;  row_3[5]  <= 16'h0842;  row_3[6]  <= 16'h0842;  row_3[7]  <= 16'h0842;
            row_3[8]  <= 16'h0846;  row_3[9]  <= 16'h083A;  row_3[10] <= 16'h0802;  row_3[11] <= 16'h0802;
            row_3[12] <= 16'h0824;  row_3[13] <= 16'h3E18;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd20: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h3C18;
            row_3[4]  <= 16'h4224;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4242;  row_3[7]  <= 16'h0242;
            row_3[8]  <= 16'h0442;  row_3[9]  <= 16'h0842;  row_3[10] <= 16'h1042;  row_3[11] <= 16'h2042;
            row_3[12] <= 16'h4224;  row_3[13] <= 16'h7E18;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd21: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h3C08;
            row_3[4]  <= 16'h4238;  row_3[5]  <= 16'h4208;  row_3[6]  <= 16'h4208;  row_3[7]  <= 16'h0208;
            row_3[8]  <= 16'h0408;  row_3[9]  <= 16'h0808;  row_3[10] <= 16'h1008;  row_3[11] <= 16'h2008;
            row_3[12] <= 16'h4208;  row_3[13] <= 16'h7E3E;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd22: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h3C3C;
            row_3[4]  <= 16'h4242;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4242;  row_3[7]  <= 16'h0202;
            row_3[8]  <= 16'h0404;  row_3[9]  <= 16'h0808;  row_3[10] <= 16'h1010;  row_3[11] <= 16'h2020;
            row_3[12] <= 16'h4242;  row_3[13] <= 16'h7E7E;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        6'd23: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h3C3C;
            row_3[4]  <= 16'h4242;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4202;  row_3[7]  <= 16'h0204;
            row_3[8]  <= 16'h0418;  row_3[9]  <= 16'h0804;  row_3[10] <= 16'h1002;  row_3[11] <= 16'h2042;
            row_3[12] <= 16'h4242;  row_3[13] <= 16'h7E3C;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
        default: begin
            row_3[0]  <= 16'h0000;  row_3[1]  <= 16'h0000;  row_3[2]  <= 16'h0000;  row_3[3]  <= 16'h1818;
            row_3[4]  <= 16'h2424;  row_3[5]  <= 16'h4242;  row_3[6]  <= 16'h4242;  row_3[7]  <= 16'h4242;
            row_3[8]  <= 16'h4242;  row_3[9]  <= 16'h4242;  row_3[10] <= 16'h4242;  row_3[11] <= 16'h4242;
            row_3[12] <= 16'h2424;  row_3[13] <= 16'h1818;  row_3[14] <= 16'h0000;  row_3[15] <= 16'h0000;
        end
    endcase
end


always @(posedge vga_clk_25 or negedge rst_n)
begin
    if(!rst_n)
        pixel_data <= WHITE;
    else begin
        
        if( ((pixel_xpos >= ROW1_X) && (pixel_xpos < ROW1_X+ROW1_H))
          && ((pixel_ypos >= ROW1_Y) && (pixel_ypos < ROW1_Y+ROW1_V)) ) begin
            if(row_1[y1_cnt][10'd159 - x1_cnt])  
                pixel_data <= RED;              
            else
                pixel_data <= WHITE;           
        end  
        
        else if( ((pixel_xpos >= ROW2_X) && (pixel_xpos < ROW2_X+ROW2_H))
               && ((pixel_ypos >= ROW2_Y) && (pixel_ypos < ROW2_Y+ROW2_V)) ) begin
                   if(row_2[y2_cnt][10'd48 - x2_cnt])  
                       pixel_data <= BLANK;              
                    else
                       pixel_data <= WHITE;           
        end 
        
        else if( ((pixel_xpos >= ROW3_X) && (pixel_xpos < ROW3_X+ROW3_H))
               && ((pixel_ypos >= ROW3_Y) && (pixel_ypos < ROW3_Y+ROW3_V)) ) begin
                   if(row_3[y3_cnt][10'd16 - x3_cnt])  
                       pixel_data <= BLANK;              
                    else
                       pixel_data <= WHITE;           
        end 
        else
            pixel_data <= WHITE;               
    end
end

endmodule 